module UARTRX #(parameter CLK_PER_BITS=1086,
                parameter IDLE=3'b000,
                parameter START=3'b001,
                parameter DATA=3'b010,
                parameter STOP=3'b011,
                 parameter CLEANUP=3'b100)
                 (input clk,input data_in,output reg[7:0] data_out,output reg dv,output reg[7:0] count,output reg[7:0] bitindex,output reg[2:0] STATE);
  
 /* parameter IDLE=3'b000;
  parameter START=3'b001;
  parameter DATA=3'b010;
  parameter STOP=3'b011;
  parameter CLEANUP=3'b100; */
  always@(posedge clk) begin
    case(STATE)
      IDLE:begin
        count<=0;
        dv<=1'b0;
        bitindex<=0;  
        if(data_in==1'b0) begin
          STATE<=START;
        end else
          STATE<=IDLE;
      end
      
      START: begin
        if(count==((CLK_PER_BITS-1)/2))begin
          if(data_in==1'b0)begin
            count<=1'b0;
          STATE<=DATA;
            
          end   
          else
            STATE<=IDLE;
        end else begin
          count<=count+1;
          STATE<=START;
        end
      end
      
      DATA: begin
     if(count<(CLK_PER_BITS)) begin
        //if(count<((CLK_PER_BITS-1)/2)) begin
        count<=count+1;
        STATE<=DATA;
     end else begin
        count<=0;
        data_out[bitindex]<=data_in;
        if (bitindex<7)
        begin
            bitindex=bitindex+1;
            STATE<=DATA;
        end else begin
            bitindex=0;
            count<=0;   
             STATE<=STOP;
             
      end
     end
      end

      
      STOP: begin
        if(count<(CLK_PER_BITS))begin
           // if(count<((CLK_PER_BITS-1)/2)) begin
            count<=count+1;
            STATE<=STOP;
        end else begin
            dv<=1'b1;
            count<=0;
        STATE<=CLEANUP;
        
      end
      end
      
      CLEANUP: begin
        dv<=1'b0;
        STATE<=IDLE;
         
      end
      
      default:
        STATE<=IDLE;
    endcase
  end
  endmodule
    
          
          
          
     
        
          
         
 
  
  